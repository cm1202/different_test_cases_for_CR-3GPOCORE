module chu_gpo
   #(parameter W = 8)  // width of output port
   (
    input  logic clk,
    input  logic reset,
    // slot interface
    input  logic cs,
    input  logic read,
    input  logic write,
    input  logic [4:0] addr,
    input  logic [31:0] wr_data,
    output logic [31:0] rd_data,
    // external port    
    output logic [W-1:0] dout
   );

   // declaration
   logic [W-1:0] buf_reg;
   logic [15:0] speed_reg;
   logic wr_en,wr_D,wr_S;

   // body
   // output buffer register
   always_ff @(posedge clk, posedge reset)
      if (reset)
         buf_reg <= 0;
      else   
         if (wr_S) begin
            speed_reg <= wr_data[15:0];
         end
      
   // decoding logic 
   assign dout[W-1:1] = 0;
   assign wr_S = cs && write && (addr == 5'b00001);
   assign rd_data =  0;
   
   blink_controller led0(
    .clk(clk),
    .rst(reset),
    .speed(speed_reg),
    .led(dout[0])
    ); 
   
   
endmodule
       



